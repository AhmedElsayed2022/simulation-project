** Profile: "SCHEMATIC1-Noninvertin OpAmp"  [ C:\USERS\EL GOHARY\ORCAD\Noninvertin OpAmp-PSpiceFiles\SCHEMATIC1\Noninvertin OpAmp.sim ] 

** Creating circuit file "Noninvertin OpAmp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\EL GOHARY\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10m 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
