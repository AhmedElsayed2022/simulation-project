** Profile: "SCHEMATIC1-Hartely oscillator"  [ C:\Users\EL GOHARY\orcad\Hartely oscillator-PSpiceFiles\HARTELY OSCILLATOR-SCHEMATIC1-Hartely oscillator.sim ] 

** Creating circuit file "HARTELY OSCILLATOR-SCHEMATIC1-Hartely oscillator.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\EL GOHARY\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 25m 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\HARTELY OSCILLATOR-SCHEMATIC1.net" 


.END
